// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 17.0.0 Build 595 04/25/2017 SJ Standard Edition
// Created on Tue Nov 14 13:28:38 2017

// synthesis message_off 10175

`timescale 1ns/1ns

module cLock (
    input reset, input clock, input C, input Enter, input Max,
    output Corr, output Err);

    enum int unsigned { corr0_err0_2=0, corr0_err1=1, corr0_err0=2, corr1_err0=3 } fstate, reg_fstate;

    always_ff @(posedge clock or posedge reset)
    begin
        if (reset) begin
            fstate <= corr0_err0;
        end
        else begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        Corr <= 1'b0;
        Err <= 1'b0;
        case (fstate)
            corr0_err0_2: begin
                if (((Enter == 1'b1) & (Max == 1'b1)))
                    reg_fstate <= corr0_err1;
                else if (((Max == 1'b0) | (Enter == 1'b0)))
                    reg_fstate <= corr0_err0_2;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= corr0_err0_2;

                Corr <= 1'b0;

                Err <= 1'b0;
            end
            corr0_err1: begin
                reg_fstate <= corr0_err1;

                Corr <= 1'b0;

                Err <= 1'b1;
            end
            corr0_err0: begin
                if ((((C == 1'b1) & (Enter == 1'b1)) & (Max == 1'b1)))
                    reg_fstate <= corr1_err0;
                else if ((((C == 1'b0) & (Enter == 1'b1)) & (Max == 1'b0)))
                    reg_fstate <= corr0_err0_2;
                else if ((((C == 1'b0) & (Enter == 1'b1)) & (Max == 1'b1)))
                    reg_fstate <= corr0_err1;
                else if (((Enter == 1'b0) | (((C == 1'b1) & (Enter == 1'b1)) & (Max == 1'b0))))
                    reg_fstate <= corr0_err0;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= corr0_err0;

                Corr <= 1'b0;

                Err <= 1'b0;
            end
            corr1_err0: begin
                reg_fstate <= corr1_err0;

                Corr <= 1'b1;

                Err <= 1'b0;
            end
            default: begin
                Corr <= 1'bx;
                Err <= 1'bx;
                $display ("Reach undefined state");
            end
        endcase
    end
endmodule // cLock
