// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 15.1.0 Build 185 10/21/2015 SJ Lite Edition
// Created on Fri Dec 08 13:06:10 2017

// synthesis message_off 10175

`timescale 1ns/1ns

module SM1 (
    input reset, input clock, input Enter, input TL,
    output R3, output R2, output R1, output R0, output Sel, output OtherEnter);

    enum int unsigned { state1=0, state2=1, state3=2, state5=3, state4=4, state6=5 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= state1;
            R3 <= 1'b0;
            R2 <= 1'b0;
            R1 <= 1'b0;
            R0 <= 1'b0;
            Sel <= 1'b0;
            OtherEnter <= 1'b0;
        end
        else begin
            R3 <= 1'b0;
            R2 <= 1'b0;
            R1 <= 1'b0;
            R0 <= 1'b0;
            Sel <= 1'b0;
            OtherEnter <= 1'b0;
            case (fstate)
                state1: begin
                    if ((Enter == 1'b1))
                        reg_fstate <= state2;
                    else if ((Enter == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    Sel <= 1'b0;

                    R1 <= 1'b1;

                    R2 <= 1'b1;

                    R0 <= 1'b1;

                    R3 <= 1'b1;

                    if ((Enter == 1'b1))
                        OtherEnter <= 1'b1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        OtherEnter <= 1'b0;
                end
                state2: begin
                    if (((TL == 1'b1) & (Enter == 1'b0)))
                        reg_fstate <= state5;
                    else if ((Enter == 1'b1))
                        reg_fstate <= state6;
                    else if (((TL == 1'b0) & (Enter == 1'b0)))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    Sel <= 1'b1;

                    R1 <= 1'b0;

                    R2 <= 1'b0;

                    R0 <= 1'b0;

                    R3 <= 1'b1;

                    if ((Enter == 1'b1))
                        OtherEnter <= 1'b1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        OtherEnter <= 1'b0;
                end
                state3: begin
                    if (((TL == 1'b1) & (Enter == 1'b0)))
                        reg_fstate <= state2;
                    else if ((Enter == 1'b1))
                        reg_fstate <= state6;
                    else if (((TL == 1'b0) & (Enter == 1'b0)))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    Sel <= 1'b1;

                    R1 <= 1'b0;

                    R2 <= 1'b0;

                    R0 <= 1'b1;

                    R3 <= 1'b0;

                    if ((Enter == 1'b1))
                        OtherEnter <= 1'b1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        OtherEnter <= 1'b0;
                end
                state5: begin
                    if ((Enter == 1'b1))
                        reg_fstate <= state6;
                    else if (((TL == 1'b1) & (Enter == 1'b0)))
                        reg_fstate <= state4;
                    else if (((TL == 1'b0) & (Enter == 1'b0)))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    Sel <= 1'b1;

                    R1 <= 1'b0;

                    R2 <= 1'b1;

                    R0 <= 1'b0;

                    R3 <= 1'b0;

                    if ((Enter == 1'b1))
                        OtherEnter <= 1'b1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        OtherEnter <= 1'b0;
                end
                state4: begin
                    if ((Enter == 1'b1))
                        reg_fstate <= state6;
                    else if (((TL == 1'b1) & (Enter == 1'b0)))
                        reg_fstate <= state3;
                    else if (((TL == 1'b0) & (Enter == 1'b0)))
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    Sel <= 1'b1;

                    R1 <= 1'b1;

                    R2 <= 1'b0;

                    R0 <= 1'b0;

                    R3 <= 1'b0;

                    if ((Enter == 1'b1))
                        OtherEnter <= 1'b1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        OtherEnter <= 1'b0;
                end
                state6: begin
                    if ((Enter == 1'b0))
                        reg_fstate <= state1;
                    else if ((Enter == 1'b1))
                        reg_fstate <= state6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state6;

                    Sel <= 1'b1;

                    R1 <= 1'b1;

                    R2 <= 1'b1;

                    R0 <= 1'b1;

                    R3 <= 1'b1;

                    OtherEnter <= 1'b0;
                end
                default: begin
                    R3 <= 1'bx;
                    R2 <= 1'bx;
                    R1 <= 1'bx;
                    R0 <= 1'bx;
                    Sel <= 1'bx;
                    OtherEnter <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM1
