// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 15.1.0 Build 185 10/21/2015 SJ Lite Edition
// Created on Fri Dec 08 12:36:54 2017

// synthesis message_off 10175

`timescale 1ns/1ns

module SM2 (
    input reset, input clock, input Enter, input Sel,
    output Pulse);

    enum int unsigned { state2=0, Columns=1, state1=2, state3=3, state4=4 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= Columns;
            Pulse <= 1'b0;
        end
        else begin
            Pulse <= 1'b0;
            case (fstate)
                state2: begin
                    if (((Sel == 1'b1) & (Enter == 1'b1)))
                        reg_fstate <= state2;
                    else if (((Sel == 1'b0) & (Enter == 1'b1)))
                        reg_fstate <= state1;
                    else if (((Enter == 1'b0) & (Sel == 1'b1)))
                        reg_fstate <= state3;
                    else if (((Sel == 1'b0) & (Enter == 1'b0)))
                        reg_fstate <= Columns;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    Pulse <= 1'b1;
                end
                Columns: begin
                    if ((Enter == 1'b0))
                        reg_fstate <= Columns;
                    else if ((Enter == 1'b1))
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Columns;

                    Pulse <= 1'b0;
                end
                state1: begin
                    if ((Enter == 1'b1))
                        reg_fstate <= state1;
                    else if ((Enter == 1'b0))
                        reg_fstate <= Columns;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    Pulse <= 1'b0;
                end
                state3: begin
                    if ((Enter == 1'b0))
                        reg_fstate <= state3;
                    else if ((Enter == 1'b1))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    Pulse <= 1'b0;
                end
                state4: begin
                    reg_fstate <= state2;

                    Pulse <= 1'b1;
                end
                default: begin
                    Pulse <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM2
